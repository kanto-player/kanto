library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sram_rom_dummy is
    port (addr : in std_logic_vector(17 downto 0);
          readdata : out std_logic_vector(15 downto 0);
          req : in std_logic;
          ack : out std_logic;
          clk : in std_logic);
end sram_rom_dummy;

architecture rtl of sram_rom_dummy is
    type state_type is (INACTIVE, RESPONDING);
    type rom_type is array(0 to 767) of std_logic_vector(15 downto 0);
    signal state : state_type := INACTIVE;
    signal rom : rom_type := (x"0000", x"04c5", x"0988", x"0e48", x"1303", x"17b7", x"1c63", x"2105", x"259b", x"2a24", x"2e9d", x"3306", x"375d", x"3ba0", x"3fce", x"43e6", x"47e5", x"4bca", x"4f95", x"5343", x"56d4", x"5a45", x"5d97", x"60c8", x"63d6", x"66c0", x"6986", x"6c26", x"6ea0", x"70f3", x"731d", x"751f", x"76f7", x"78a4", x"7a27", x"7b7e", x"7ca9", x"7da8", x"7e7a", x"7f1f", x"7f97", x"7fe2", x"7fff", x"7fef", x"7fb1", x"7f45", x"7ead", x"7de7", x"7cf5", x"7bd6", x"7a8b", x"7914", x"7773", x"75a7", x"73b1", x"7192", x"6f4b", x"6cdb", x"6a46", x"678a", x"64aa", x"61a6", x"5e7f", x"5b36", x"57cd", x"5445", x"509f", x"4cdc", x"48fe", x"4506", x"40f5", x"3ccd", x"3890", x"343e", x"2fda", x"2b65", x"26e0", x"224e", x"1db0", x"1906", x"1454", x"0f9b", x"0adc", x"061a", x"0155", x"fc90", x"f7cc", x"f30b", x"ee4e", x"e998", x"e4ea", x"e045", x"dbac", x"d71f", x"d2a1", x"ce33", x"c9d7", x"c58f", x"c15b", x"bd3d", x"b936", x"b54a", x"b177", x"adc1", x"aa28", x"a6ae", x"a353", x"a019", x"9d01", x"9a0d", x"973d", x"9492", x"920d", x"8faf", x"8d79", x"8b6c", x"8989", x"87d0", x"8641", x"84de", x"83a6", x"829b", x"81bc", x"810a", x"8086", x"802e", x"8004", x"8008", x"803a", x"8098", x"8124", x"81dd", x"82c3", x"83d6", x"8514", x"867e", x"8814", x"89d4", x"8bbf", x"8dd2", x"900f", x"9273", x"94fd", x"97af", x"9a85", x"9d7f", x"a09c", x"a3dc", x"a73c", x"aabb", x"ae59", x"b214", x"b5eb", x"b9dc", x"bde6", x"c207", x"c63f", x"ca8b", x"ceea", x"d35a", x"d7db", x"dc6a", x"e105", x"e5ab", x"ea5b", x"ef13", x"f3d0", x"f892", x"fd56", x"021b", x"06df", x"0ba1", x"1060", x"1518", x"19c8", x"1e70", x"230d", x"279d", x"2c1f", x"3092", x"34f3", x"3941", x"3d7b", x"419f", x"45ac", x"49a0", x"4d7a", x"5138", x"54da", x"585d", x"5bc1", x"5f04", x"6225", x"6523", x"67fe", x"6ab4", x"6d43", x"6fac", x"71ed", x"7405", x"75f4", x"77b9", x"7954", x"7ac4", x"7c07", x"7d1f", x"7e0a", x"7ec9", x"7f5a", x"7fbe", x"7ff4", x"7ffe", x"7fd9", x"7f87", x"7f08", x"7e5b", x"7d82", x"7c7c", x"7b49", x"79eb", x"7861", x"76ad", x"74cf", x"72c6", x"7095", x"6e3c", x"6bbc", x"6916", x"664a", x"6359", x"6046", x"5d10", x"59b9", x"5642", x"52ac", x"4ef9", x"4b2b", x"4740", x"433e", x"3f22", x"3af1", x"36aa", x"3251", x"2de5", x"2969", x"24de", x"2046", x"1ba2", x"16f5", x"1240", x"0d83", x"08c3", x"03ff", x"ff3b", x"fa76", x"f5b3", x"f0f3", x"ec39", x"e786", x"e2dc", x"de3c", x"d9a8", x"d522", x"d0ab", x"cc45", x"c7f1", x"c3b1", x"bf87", x"bb73", x"b778", x"b397", x"afd1", x"ac27", x"a89b", x"a52f", x"a1e2", x"9eb7", x"9baf", x"98ca", x"960a", x"9370", x"90fc", x"8eb0", x"8c8d", x"8a92", x"88c1", x"871a", x"859f", x"844f", x"832b", x"8233", x"8168", x"80ca", x"805a", x"8016", x"8000", x"8018", x"805e", x"80d0", x"8170", x"823d", x"8337", x"845d", x"85af", x"872c", x"88d5", x"8aa8", x"8ca4", x"8eca", x"9118", x"938d", x"9629", x"98eb", x"9bd1", x"9edb", x"a207", x"a555", x"a8c3", x"ac50", x"affb", x"b3c3", x"b7a5", x"bba1", x"bfb6", x"c3e1", x"c822", x"cc76", x"d0dd", x"d555", x"d9dc", x"de71", x"e311", x"e7bc", x"ec6f", x"f129", x"f5e9", x"faac", x"ff71", x"0435", x"08f9", x"0dba", x"1276", x"172b", x"1bd8", x"207a", x"2512", x"299c", x"2e18", x"3283", x"36dc", x"3b21", x"3f52", x"436c", x"476e", x"4b56", x"4f24", x"52d6", x"566a", x"59e0", x"5d35", x"606a", x"637c", x"666a", x"6935", x"6bd9", x"6e58", x"70af", x"72de", x"74e5", x"76c1", x"7874", x"79fc", x"7b58", x"7c88", x"7d8c", x"7e64", x"7f0e", x"7f8c", x"7fdb", x"7ffe", x"7ff3", x"7fba", x"7f54", x"7ec1", x"7e01", x"7d13", x"7bfa", x"7ab4", x"7943", x"77a6", x"75df", x"73ee", x"71d4", x"6f91", x"6d26", x"6a95", x"67de", x"6502", x"6202", x"5edf", x"5b9b", x"5835", x"54b1", x"510e", x"4d4e", x"4973", x"457e", x"4170", x"3d4b", x"3910", x"34c1", x"305f", x"2bec", x"2769", x"22d8", x"1e3b", x"1993", x"14e2", x"1029", x"0b6b", x"06a9", x"01e4", x"fd20", x"f85b", x"f39a", x"eedc", x"ea25", x"e576", x"e0d0", x"dc35", x"d7a7", x"d327", x"ceb8", x"ca59", x"c60e", x"c1d7", x"bdb7", x"b9ae", x"b5be", x"b1e9", x"ae2f", x"aa92", x"a714", x"a3b6", x"a078", x"9d5c", x"9a64", x"978f", x"94e0", x"9257", x"8ff4", x"8dba", x"8ba8", x"89bf", x"8801", x"866d", x"8505", x"83c8", x"82b8", x"81d4", x"811d", x"8093", x"8036", x"8007", x"8005", x"8031", x"808a", x"8111", x"81c5", x"82a6", x"83b3", x"84ec", x"8652", x"87e2", x"899e", x"8b83", x"8d92", x"8fc9", x"9229", x"94af", x"975c", x"9a2e", x"9d24", x"a03d", x"a379", x"a6d5", x"aa51", x"adeb", x"b1a3", x"b576", x"b964", x"bd6b", x"c18a", x"c5bf", x"ca09", x"ce66", x"d2d4", x"d753", x"dbe0", x"e07a", x"e51f", x"e9ce", x"ee84", x"f341", x"f803", x"fcc7", x"018b", x"0650", x"0b13", x"0fd1", x"148a", x"193c", x"1de5", x"2283", x"2715", x"2b99", x"300d", x"3470", x"38c1", x"3cfd", x"4124", x"4534", x"492b", x"4d08", x"50c9", x"546e", x"57f5", x"5b5d", x"5ea4", x"61c9", x"64cc", x"67aa", x"6a64", x"6cf8", x"6f65", x"71ab", x"73c8", x"75bc", x"7787", x"7926", x"7a9b", x"7be4", x"7d00", x"7df1", x"7eb5", x"7f4b", x"7fb4", x"7ff0", x"7fff", x"7fe0", x"7f93", x"7f19", x"7e72", x"7d9d", x"7c9d", x"7b6f", x"7a16", x"7892", x"76e2", x"7509", x"7305", x"70d9", x"6e85", x"6c09", x"6967", x"66a0", x"63b3", x"60a4", x"5d72", x"5a1f", x"56ac", x"5319", x"4f6a", x"4b9e", x"47b7", x"43b7", x"3f9f", x"3b70", x"372c", x"32d4", x"2e6a", x"29f0", x"2567", x"20d0", x"1c2e", x"1782", x"12cd", x"0e12", x"0952", x"048e", x"ffca", x"fb05", x"f641", x"f182", x"ecc7", x"e813", x"e367", x"dec6", x"da31", x"d5a9", x"d130", x"ccc8", x"c872", x"c42f", x"c002", x"bbec", x"b7ee", x"b40a", x"b040", x"ac93", x"a904", x"a594", x"a244", x"9f15", x"9c08", x"991f", x"965b", x"93bc", x"9144", x"8ef3", x"8ccb", x"8acb", x"88f5", x"874a", x"85c9", x"8474", x"834b", x"824e", x"817e", x"80da", x"8064", x"801c", x"8001", x"8013", x"8053", x"80c1", x"815b", x"8223", x"8317", x"8438", x"8585", x"86fd", x"88a1", x"8a6f", x"8c66", x"8e87", x"90d1", x"9341", x"95d9", x"9896", x"9b78", x"9e7e", x"a1a6", x"a4f0", x"a85b", x"abe4", x"af8c", x"b350", x"b72f", x"bb28", x"bf3a", x"c363", x"c7a1", x"cbf3", x"d058", x"d4ce", x"d953", x"dde6", x"e286", x"e72f", x"ebe2", x"f09b", x"f55a", x"fa1d", x"fee2", x"03a6", x"086a", x"0d2b", x"11e8", x"169e", x"1b4c", x"1ff0", x"2489", x"2915", x"2d92", x"31ff", x"365a", x"3aa2", x"3ed5", x"42f2", x"46f7", x"4ae2", x"4eb4", x"5269", x"5600", x"597a", x"5cd3", x"600b", x"6321", x"6614", x"68e3", x"6b8c", x"6e0f", x"706b", x"729f", x"74aa", x"768c", x"7843", x"79d0", x"7b31", x"7c67", x"7d70", x"7e4d", x"7efd", x"7f7f", x"7fd5", x"7ffc", x"7ff7", x"7fc3", x"7f63", x"7ed5", x"7e1a", x"7d32", x"7c1d", x"7add", x"7970", x"77d9", x"7617", x"742a", x"7215", x"6fd7", x"6d71", x"6ae4", x"6832", x"655a", x"625e", x"5f3f", x"5bfe", x"589d", x"551c", x"517d", x"4dc0", x"49e9", x"45f6", x"41eb", x"3dc9", x"3991", x"3544", x"30e4", x"2c72", x"27f1", x"2362", x"1ec6", x"1a1f", x"156f", x"10b7", x"0bfa", x"0738", x"0273", x"fdaf", x"f8ea", x"f428", x"ef6a", x"eab3", x"e602", x"e15b", x"dcbf", x"d82f");
    signal intern_addr : unsigned(17 downto 0);
begin
    intern_addr <= unsigned(addr);
    process (clk)
    begin
        if rising_edge(clk) then
            case state is
                when INACTIVE =>
                    if req = '1' then
                        state <= RESPONDING;
                    end if;
                when RESPONDING =>
                    if req = '0' then
                        state <= INACTIVE;
                    end if;
            end case;
        end if;
    end process;
    
    readdata <= rom(to_integer(intern_addr)) 
                    when state = responding else x"0000";
    ack <= '1' when state = RESPONDING else '0';
end rtl;
