// de2_vga_text_buffer_0.v

// Generated using ACDS version 12.1 177 at 2013.05.13.12:49:07

`timescale 1 ps / 1 ps
module de2_vga_text_buffer_0 (
		input  wire         vga_read,         //         vga.read
		input  wire         vga_write,        //            .write
		input  wire         vga_chipselect,   //            .chipselect
		input  wire [9:0]   vga_address,      //            .address
		output wire [127:0] vga_readdata,     //            .readdata
		input  wire [127:0] vga_writedata,    //            .writedata
		input  wire         vga_clk,          //  clock_sink.clk
		input  wire         vga_reset,        //  reset_sink.reset
		output wire         display_pixel_on  // conduit_end.export
	);

	de2_vga_text_buffer de2_vga_text_buffer_0_inst (
		.vga_read         (vga_read),         //         vga.read
		.vga_write        (vga_write),        //            .write
		.vga_chipselect   (vga_chipselect),   //            .chipselect
		.vga_address      (vga_address),      //            .address
		.vga_readdata     (vga_readdata),     //            .readdata
		.vga_writedata    (vga_writedata),    //            .writedata
		.vga_clk          (vga_clk),          //  clock_sink.clk
		.vga_reset        (vga_reset),        //  reset_sink.reset
		.display_pixel_on (display_pixel_on)  // conduit_end.export
	);

endmodule
