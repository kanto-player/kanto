// ps2.v

// Generated using ACDS version 12.1 177 at 2013.05.13.07:12:33

`timescale 1 ps / 1 ps
module ps2 (
		input  wire [2:0] avs_s1_address,    // avalon_slave_0.address
		input  wire       avs_s1_read,       //               .read
		input  wire       avs_s1_chipselect, //               .chipselect
		output wire [7:0] avs_s1_readdata,   //               .readdata
		input  wire       PS2_Clk,           //    conduit_end.export
		input  wire       PS2_Data,          //               .export
		input  wire       avs_s1_clk,        //     clock_sink.clk
		input  wire       avs_s1_reset       //     reset_sink.reset
	);

	de2_ps2 ps2_inst (
		.avs_s1_address    (avs_s1_address),    // avalon_slave_0.address
		.avs_s1_read       (avs_s1_read),       //               .read
		.avs_s1_chipselect (avs_s1_chipselect), //               .chipselect
		.avs_s1_readdata   (avs_s1_readdata),   //               .readdata
		.PS2_Clk           (PS2_Clk),           //    conduit_end.export
		.PS2_Data          (PS2_Data),          //               .export
		.avs_s1_clk        (avs_s1_clk),        //     clock_sink.clk
		.avs_s1_reset      (avs_s1_reset)       //     reset_sink.reset
	);

endmodule
